// Created: February 22, 2025
// Author - Aditya Vikram Singh, Shiva Shankar B

module proElement(
	input w [31:0], //weights
	input x [31:0], // input
	input b [31:0], // base

	input count [9:0], //counter for operation

	input head, //header
	input clock,

	output pe_out [31:0], // output of processing element
	output done_flag //flag when operations are done
);






endmodule

module soft_max(
    
);
endmodule